library verilog;
use verilog.vl_types.all;
entity TestBench1 is
end TestBench1;
