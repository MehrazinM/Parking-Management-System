library verilog;
use verilog.vl_types.all;
entity TestBench2 is
end TestBench2;
