library verilog;
use verilog.vl_types.all;
entity TestBench3 is
end TestBench3;
